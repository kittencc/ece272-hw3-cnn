// connects simple_read_FSM, read_addr_gen, read_bank_counter modules
// relays control signals between the read_FSM and the main_FSM
// Author: Cheryl (Yingqiu) Cao
// Date: 2022-01-2

module simple_read_controller
# (
  parameter CONFIG_WIDTH = 32,
  parameter BANK_ADDR_WIDTH = 32,
  parameter COUNTER_WID = 8,             // needs to be large enough to save IC1*IX0*IY0
  parameter OY1_OX1 = 4*4       // used for the write_bank_counter

)
(
  input logic clk,
  input logic rst_n,

  // for read_addr_gen
  input logic [CONFIG_WIDTH - 1 : 0] config_data,
 
  // for the read FSM
  input logic start_new_read_bank,
  output logic read_bank_ready_to_switch,
  output logic [COUNTER_WID - 1 : 0] read_bank_count,

  // to read from the double buffer
  output logic ren,
  output logic [BANK_ADDR_WIDTH - 1 : 0] raddr    // read addr generated by the module

);


// local signal begin
// for read_addr_gen
logic addr_enable;        // en signal
logic config_enable;
logic reading_last_data;

// for the read FSM
logic one_read_bank_done;
// local signal end


assign ren = addr_enable;        // addr gen is synced with ren of the double buffer

// connect read_bank_counter 
//  counts from 0 to MAX_COUNT - 1;
counter  
#(
  .MAX_COUNT(OY1_OX1+1),
  .COUNTER_WID(COUNTER_WID)
)
read_bank_counter_inst
(
  .clk(clk),
  .rst_n(rst_n),
  .en(one_read_bank_done),
  .count(read_bank_count)
);



// connect simple_read_FSM module
simple_read_FSM read_FSM_inst
(
  .clk(clk),
  .rst_n(rst_n),
  .start_new_read_bank(start_new_read_bank),
  .reading_last_data(reading_last_data),   
  .config_enable(config_enable),            // for the addr gen module
  .addr_enable(addr_enable),              // en signal for the addr gen module
  .one_read_bank_done(one_read_bank_done),
  .read_bank_ready_to_switch(read_bank_ready_to_switch)
);





// connect read_addr_gen inst
// in this particular tb, we are using the same read order as write
input_write_addr_gen 
#( 
  .CONFIG_WIDTH(CONFIG_WIDTH),
  .BANK_ADDR_WIDTH(BANK_ADDR_WIDTH)
)
input_read_addr_gen_inst
(
  .clk(clk),
  .rst_n(rst_n),
  .addr_enable(addr_enable),
  .config_enable(config_enable),
  .config_data(config_data),
  .addr(raddr),
  .writing_last_data(reading_last_data)
);



endmodule
